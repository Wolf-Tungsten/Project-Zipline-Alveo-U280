/*************************************************************************
*
* Copyright � Microsoft Corporation. All rights reserved.
* Copyright � Broadcom Inc. All rights reserved.
* Licensed under the MIT License.
*
*************************************************************************/



`ifndef __CR_SU_VH
`define __CR_SU_VH


`include "cr_su_regs.vh"
`include "cr_su_regsPKG.svp"
`include "cr_su_regfilePKG.svp"
`include "cr_suPKG.svp"

`define MAX(a,b) \
    (((a)>(b))?(a):(b))
`define MIN(a,b) \
    (((a)<(b))?(a):(b))
`define LOG_VEC(a) `MAX(0, ($clog2(a)-1)):0


`endif 



    
